module main

fn print_header(s string) {
	println(s)
	println(`=`.repeat(s.len))
}
